LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_UNSIGNED.ALL;

ENTITY CLK_CTROL2 IS
  PORT(CLK_IN:IN STD_LOGIC;
       START2:IN STD_LOGIC;
		 CLK:OUT STD_LOGIC);
END CLK_CTROL2;

ARCHITECTURE ART OF CLK_CTROL2 IS
BEGIN

PROCESS(CLK_IN)IS
  BEGIN
  IF START2='1' THEN
    CLK<=CLK_IN;
  ELSE
    CLK<='0';
  END IF;
END PROCESS;
END ART;
