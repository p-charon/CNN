LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;

ENTITY REG_B IS
PORT(
     start4:IN STD_LOGIC;
	  Y:IN STD_LOGIC_VECTOR(10 DOWNTO 0);
	  Q:BUFFER STD_LOGIC_VECTOR(10 DOWNTO 0));
END ENTITY;
ARCHITECTURE ART OF REG_B IS
SIGNAL CNT:STD_LOGIC_VECTOR(10 DOWNTO 0);
BEGIN
PROCESS(Y)IS
BEGIN
  CNT<=Y;
 IF (start4='1') THEN
 Q<=CNT;
 ELSE NULL;
 END IF;
 END PROCESS;
 END ARCHITECTURE ART;