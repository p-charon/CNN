LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_SIGNED.ALL;

ENTITY SULE IS
PORT(CLK:IN STD_LOGIC;
     Q1:IN STD_LOGIC_VECTOR(10 DOWNTO 0); 
	  Y:BUFFER STD_LOGIC_VECTOR(10 DOWNTO 0));
END ENTITY;
ARCHITECTURE ART OF SULE IS
BEGIN
PROCESS(Q1,CLK)IS
BEGIN
IF CLK'EVENT AND CLK='1' THEN
IF (Q1>"00000000000") THEN
Y<=Q1;
ELSE
Y<="00000000000";
 END IF;
 END IF;
 END PROCESS;
END ARCHITECTURE ART;