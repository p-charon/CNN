LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;
USE IEEE.STD_LOGIC_UNSIGNED.ALL;

ENTITY CARRAY3232 IS
GENERIC( W1:INTEGER:=11;   --样本位宽
			W3:INTEGER:=784;  --样本数组长度
			W4:INTEGER:=196); --输出数组长度

 PORT(CLK:IN STD_LOGIC;
		START2:IN STD_LOGIC;
		OVER2:OUT STD_LOGIC;
      OUTA:OUT STD_LOGIC_VECTOR(W1-1 DOWNTO 0);
		OUTB:OUT STD_LOGIC_VECTOR(W1-1 DOWNTO 0);
		OUTC:OUT STD_LOGIC_VECTOR(W1-1 DOWNTO 0);
		OUTD:OUT STD_LOGIC_VECTOR(W1-1 DOWNTO 0);
		OUTE:OUT STD_LOGIC_VECTOR(W1-1 DOWNTO 0);
		SAMENTER:IN STD_LOGIC_VECTOR(W1-1 DOWNTO 0));--样本输入
END ENTITY;

ARCHITECTURE ART OF CARRAY3232 IS
 SUBTYPE N1 IS STD_LOGIC_VECTOR(W1-1 DOWNTO 0);  --样本数组宽度
 TYPE ARRAY_N1 IS ARRAY(0 TO W3-1) OF N1;  --样本数组长度
 TYPE ARRAY_N3 IS ARRAY(0 TO W4-1) OF N1;	 --输出数组长度

 SIGNAL SAMARRAY:ARRAY_N1;		 --样本矩阵
 SIGNAL OUTARRAY:ARRAY_N3;		--输出矩阵
 SIGNAL OUTARRAY1:ARRAY_N3;

 SIGNAL A:INTEGER RANGE 0 TO W3;
 SIGNAL E:INTEGER RANGE 0 TO W4;
 SIGNAL X:INTEGER RANGE 0 TO W4;
 SIGNAL N:INTEGER RANGE 0 TO 14;
 SIGNAL Y:INTEGER RANGE 0 TO 13;
 SIGNAL COUNT:INTEGER RANGE 0 TO 4;
 SIGNAL J,C,D:STD_LOGIC:='0';
 
 BEGIN

 LOAD:PROCESS(CLK,SAMENTER,A) IS
  BEGIN 
  IF START2='1' THEN
  IF CLK'EVENT AND CLK='1' THEN
   IF A<W3 THEN	
      A<=A+1;
		C<='0';
	ELSE
	   C<='1';
	--	A<=0;
  END IF;
  SAMARRAY(A)<=SAMENTER;
  END IF;
  END IF;
END PROCESS;
 
 JISUAN:PROCESS(SAMARRAY,N,CLK) IS
  BEGIN
  IF C='1' THEN 
  IF CLK'EVENT AND CLK='1' THEN
	 FOR Y IN 0 TO 13 LOOP
	 OUTARRAY(14*N+Y)<=SAMARRAY(56*N+2*Y)+SAMARRAY(56*N+2*Y+1)+SAMARRAY(56*N+2*Y+28)+SAMARRAY(24*N+2*Y+29);
	 END LOOP;
	 N<=N+1;
	END IF;
  END IF;
  
  IF N=14 THEN
     D<='1';
  ELSE 
     D<='0';
  END IF;
  END PROCESS;
  
  CUNCHU:PROCESS(CLK,D)
  BEGIN
  	IF D='1' THEN
   IF CLK'EVENT AND CLK='1' THEN
	  IF CONV_INTEGER(OUTARRAY(E)(W1-1)&"00"&OUTARRAY(E)(W1-2 DOWNTO 2))>0 THEN
	     OUTARRAY1(E)<=OUTARRAY(E)(W1-1)&"00"&OUTARRAY(E)(W1-2 DOWNTO 2);
		ELSE
		  OUTARRAY1(E)<="00000000000";
		END IF;
		E<=E+1;
		END IF;
	END IF;
	END PROCESS;
	
	PROCESS(J) IS
	BEGIN
		IF E>196 THEN
		J<='1';
	ELSE
		J<='0';
	END IF;
	END PROCESS;
	
	PROCESS(CLK,X,COUNT) IS
	BEGIN
	IF J='1' THEN
		OVER2<='1';
	IF CLK'EVENT AND CLK='1' THEN
	 IF COUNT<5 THEN
		COUNT<=COUNT+1;
		X<=X+1;
		OUTA<=OUTARRAY1(X+14*0);
		OUTB<=OUTARRAY1(X+14*1);
		OUTC<=OUTARRAY1(X+14*2);
		OUTD<=OUTARRAY1(X+14*3);
		OUTE<=OUTARRAY1(X+14*4);
	 ELSIF  (x REM 14)/=0 THEN
				X<=X-3;
				COUNT<=1;
				OUTA<=OUTARRAY1(X-4+14*0);
				OUTB<=OUTARRAY1(X-4+14*1);
				OUTC<=OUTARRAY1(X-4+14*2);
				OUTD<=OUTARRAY1(X-4+14*3);
				OUTE<=OUTARRAY1(X-4+14*4);
		ELSE
				OUTA<=OUTARRAY1(X+14*0);
				OUTB<=OUTARRAY1(X+14*1);
				OUTC<=OUTARRAY1(X+14*2);
				OUTD<=OUTARRAY1(X+14*3);
				OUTE<=OUTARRAY1(X+14*4);
				X<=X+1;
				COUNT<=1;
		END IF;
		
	IF X>140 THEN
		X<=140;
		OUTA<="ZZZZZZZZZZZ";
		OUTB<="ZZZZZZZZZZZ";
		OUTC<="ZZZZZZZZZZZ";
		OUTD<="ZZZZZZZZZZZ";
		OUTE<="ZZZZZZZZZZZ";
	END IF;

	IF X=140 THEN
		OUTA<="ZZZZZZZZZZZ";
		OUTB<="ZZZZZZZZZZZ";
		OUTC<="ZZZZZZZZZZZ";
		OUTD<="ZZZZZZZZZZZ";
		OUTE<="ZZZZZZZZZZZ";
	END IF;
		
	END IF;
	END IF;
  END PROCESS;
END ARCHITECTURE;