LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_UNSIGNED.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

ENTITY INTIAL IS
  GENERIC (W1 : INTEGER := 9; 
           W2 : INTEGER := 1024);
  PORT(DATAIN:IN STD_LOGIC_VECTOR(W1-1 DOWNTO 0);
       CLK:IN STD_LOGIC;
		 RES:IN STD_LOGIC;
		 start:IN STD_LOGIC;
		 over1:OUT STD_LOGIC;
		 TEXTA:OUT STD_LOGIC_VECTOR(W1-1 DOWNTO 0);
		 TEXTB:OUT STD_LOGIC_VECTOR(W1-1 DOWNTO 0);
		 OUTA:OUT STD_LOGIC_VECTOR(W1-1 DOWNTO 0);
		 OUTB:OUT STD_LOGIC_VECTOR(W1-1 DOWNTO 0);
		 OUTC:OUT STD_LOGIC_VECTOR(W1-1 DOWNTO 0);
		 OUTD:OUT STD_LOGIC_VECTOR(W1-1 DOWNTO 0);
		 OUTE:OUT STD_LOGIC_VECTOR(W1-1 DOWNTO 0));
END INTIAL;

ARCHITECTURE ART OF INTIAL IS

  SUBTYPE N1BIT IS STD_LOGIC_VECTOR(W1-1 DOWNTO 0);
  TYPE DATA_N1BIT IS ARRAY (0 TO W2-1) OF N1BIT;
  SIGNAL  C  :  DATA_N1BIT; 
  SIGNAL  TEMP1:INTEGER RANGE 0 TO W2;
  SIGNAL  TEMP2:INTEGER RANGE 0 TO W2;
  SIGNAL  X,X2:INTEGER RANGE 0 TO 1025;
  SIGNAL  CONTROL:STD_LOGIC;
  SIGNAL  COUNT2:INTEGER RANGE 1 TO 5;
  SIGNAL  COUNT:INTEGER RANGE 1 TO 28;
    BEGIN
  
  LOAD:PROCESS(CLK,RES)
  BEGIN
    IF start='1' THEN
	  IF RES='0' THEN
	    FOR I IN 0 TO 1023 LOOP
		 C(I)<=(OTHERS=>'0');
		 END LOOP;
		 
		 ELSIF CLK'EVENT AND CLK='1' THEN
		 IF COUNT<28 THEN
		   COUNT<=COUNT+1;
		   X<=X+1;
		   C(34+X)<=DATAIN;
			TEMP1<=34+X;
			
		   ELSIF COUNT=28 THEN
			COUNT<=1;
			X<=X+5;
			C(34+X)<=DATAIN;
			TEMP1<=34+X;
		 END IF;
		END IF;
     END IF;
	  
	  
	 IF CLK'EVENT AND CLK='1' THEN
		IF X>=957 THEN
		  CONTROL<='1';
		ELSE 
		  CONTROL<='0';
		END IF;
	  END IF;
	  
   END PROCESS;
  
   DATAPUT:PROCESS(CLK)
	  BEGIN
	  IF CLK'EVENT AND CLK='1' THEN
	    IF CONTROL='1' THEN
	     IF COUNT2<5 THEN
			 COUNT2<=COUNT2+1;
			 OUTA<=C(X2+32*0);
			 OUTB<=C(X2+32*1);
			 OUTC<=C(X2+32*2);
			 OUTD<=C(X2+32*3);
			 OUTE<=C(X2+32*4);
			 TEMP2<=X2;
			 X2<=X2+1;
		    ELSIF  ((X2+1) REM 32)/=0 THEN
				 COUNT2<=1;
				 OUTA<=C(X2+32*0);
				 OUTB<=C(X2+32*1);
				 OUTC<=C(X2+32*2);
				 OUTD<=C(X2+32*3);
				 OUTE<=C(X2+32*4);
				 TEMP2<=X2;
				 X2<=X2+1;
			  ELSE
				 OUTA<=C(X2+32*0);
				 OUTB<=C(X2+32*1);
				 OUTC<=C(X2+32*2);
				 OUTD<=C(X2+32*3);
				 OUTE<=C(X2+32*4);
				 TEMP2<=X2;
				 X2<=X2-3;
				 COUNT2<=1;
		    END IF;

		  END IF;
	  END IF;
	END PROCESS;
  over1<=CONTROL;
  TEXTA<=CONV_STD_LOGIC_VECTOR(TEMP1,W1);
  TEXTB<=CONV_STD_LOGIC_VECTOR(TEMP2,W1);
END ART;